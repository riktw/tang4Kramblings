-- megafunction wizard: %RAM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: InternalRam4K.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity InternalRam4K is
  
  port(
        address		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
        clock		: IN STD_LOGIC  := '1';
        data		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        wren		: IN STD_LOGIC ;
        q		    : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
    );
end InternalRam4K;

architecture arch of InternalRam4K is
 type ram_type is array (2**10 downto 0) of std_logic_vector (7 downto 0);
 signal ram_single_port : ram_type;
begin
  process(clock)
  begin 
    if (clock'event and clock='1') then
      if (wren='1') then -- write data to address 'addr'
        --convert 'addr' type to integer from std_logic_vector
        ram_single_port(to_integer(unsigned(address))) <= data;
      end if;
  end if;
  end process;

  -- read data from address 'addr'
  -- convert 'addr' type to integer from std_logic_vector
  q<=ram_single_port(to_integer(unsigned(address)));
end arch;
