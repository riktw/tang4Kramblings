-- megafunction wizard: %ROM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: M6502_BASIC_ROM.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;
use ieee.std_logic_misc.ALL;
use std.textio.all;
use ieee.std_logic_textio.all;


ENTITY M6502_BASIC_ROM IS
	PORT
	(
		address		: IN STD_LOGIC_VECTOR (12 DOWNTO 0);
		clock		: IN STD_LOGIC  := '1';
		q		    : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END M6502_BASIC_ROM;


ARCHITECTURE SYN OF m6502_basic_rom IS

    type rom_array is array((2**12)-1 downto 0)
        of std_logic_vector(7 downto 0);
     
    impure function rom_init(filename : string) return rom_array is
      file rom_file : text open read_mode is filename;
      variable rom_line : line;
      variable rom_value : bit_vector(7 downto 0);
      variable temp : rom_array;
    begin
      for rom_index in 0 to (2**12)-1 loop
        readline(rom_file, rom_line);
        hread(rom_line, temp(rom_index));
      end loop;
      return temp;
    end function;
     
    signal ram : rom_array := rom_init(filename => "/mnt/80217a00-9155-4626-a8d5-81d9da63b1e8/Git/TangNano-4K-example/multicomp/6502/src/fw.hex");
    signal addr_reg : natural range 0 to 2**12;

begin

    process(clock)
	begin
        addr_reg <= to_integer(unsigned(address));
    end process;

    q <= ram(addr_reg);

END SYN;

