--Copyright (C)2014-2021 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--GOWIN Version: V1.9.8
--Part Number: GW1NSR-LV4CQN48PC7/I6
--Device: GW1NSR-4C
--Created Time: Sun Sep 12 19:16:34 2021

library IEEE;
use IEEE.std_logic_1164.all;

entity basicRom is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(12 downto 0)
    );
end basicRom;

architecture Behavioral of basicRom is

    signal prom_inst_0_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(29 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(29 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 9;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(1 downto 0) <= prom_inst_0_DO_o(1 downto 0) ;
    prom_inst_0_dout_w(29 downto 0) <= prom_inst_0_DO_o(31 downto 2) ;
    prom_inst_1_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(3 downto 2) <= prom_inst_1_DO_o(1 downto 0) ;
    prom_inst_1_dout_w(29 downto 0) <= prom_inst_1_DO_o(31 downto 2) ;
    prom_inst_2_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(5 downto 4) <= prom_inst_2_DO_o(1 downto 0) ;
    prom_inst_2_dout_w(29 downto 0) <= prom_inst_2_DO_o(31 downto 2) ;
    prom_inst_3_AD_i <= ad(12 downto 0) & gw_gnd;
    dout(7 downto 6) <= prom_inst_3_DO_o(1 downto 0) ;
    prom_inst_3_dout_w(29 downto 0) <= prom_inst_3_DO_o(31 downto 2) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"EA460278D7349FCC8FD0C210FCF5C8ED2D2C0B0820DDC1AEBE9B9F88C606BB59",
            INIT_RAM_01 => X"40CEB093694CD0BC987C919C705C1ACCD6A469FDB3699B3C41650494406B8913",
            INIT_RAM_02 => X"C4130ED7BE3EBA0140D82423F462393521927FC1F0A9FC6ADE49BC6B26E7133A",
            INIT_RAM_03 => X"4180544EC952702DD16640DB0084B19DC745DD6605155008D6A49F9090BA49B3",
            INIT_RAM_04 => X"F0C4927300312441151113002211522008042722D02214020849536226E19406",
            INIT_RAM_05 => X"4C0159D8585CD88A90D52B14230D92D1D1DDD2491D5D99402138F18E20B8000E",
            INIT_RAM_06 => X"4D0D0C414541C1C50DE080102122594195094314093150858530093440D0D710",
            INIT_RAM_07 => X"614240249085C18044110B840801010D0D0009181100E01D10376AAAAAAB4220",
            INIT_RAM_08 => X"5853046765545050324A4809150C0990C9E94A53641018060D1B902401011810",
            INIT_RAM_09 => X"210264A4024490495D89500F00010208F104201D9DD505118991518A80D850D8",
            INIT_RAM_0A => X"D04113438A0429645345141301120102CCB4000D08336A4A4090746244DC1632",
            INIT_RAM_0B => X"1870028DD074DD20D8012734036036414D07CE2402248F1078854D55D1920F14",
            INIT_RAM_0C => X"8068208E00D850DDA302B209308914214343403504D00D121540004148074C11",
            INIT_RAM_0D => X"13413400A282C194DD4047756608A5030B432474F1890804D04D068D80833080",
            INIT_RAM_0E => X"7772988207C0280390404E1C9308CD107C1412244C900434B7840388A0A37438",
            INIT_RAM_0F => X"841C902404C9CD9400C8593326630CB22437CD0D33402A17569A65555A694156",
            INIT_RAM_10 => X"48A8841062124495AC080080336490218CC923407370730820D9364D90B32406",
            INIT_RAM_11 => X"85C936AB8280CD9C100341100C5045880A820402202C4980485F005D09040206",
            INIT_RAM_12 => X"0C003983222080E86850D0D321A443BC00CB08D6247023CDD32480D0D321400D",
            INIT_RAM_13 => X"32A1544CF2D9345D134A88E1CD0080D85850D030708C0C634F001043441D9C9D",
            INIT_RAM_14 => X"6755C44B84C000D146F138008020205034CC0024931E8C6C91BB46070C81C508",
            INIT_RAM_15 => X"64CD0D00EA00D4DD597372423470A1480B8A3A8243330092801048AD98177511",
            INIT_RAM_16 => X"4D8483040C101149378091940A1020DE03405109CDCE28EAE0CB10F080090597",
            INIT_RAM_17 => X"0334041164E0CC523274D93754C0C5F081043727340427143300D10447491413",
            INIT_RAM_18 => X"4515D53C15DD595100C804DF6790D0820E0893628D24E01008BC13B24CD0128A",
            INIT_RAM_19 => X"80210B4F3636868EC55030B20C1D20501286A2161868ED112C03447772CD1756",
            INIT_RAM_1A => X"0535140499049042761422780B546CC1508086DDC185300B14403880C508DA20",
            INIT_RAM_1B => X"50450640000411325652144C9264924906449D085105C41124C90DC985012724",
            INIT_RAM_1C => X"820B364A49224634904C01DA96934F1204815D6645466013470D0400D2440C13",
            INIT_RAM_1D => X"39B0448E10DB20C18545064DAC26241250081E9016449DA2D06C630C9056326A",
            INIT_RAM_1E => X"84764994149514648AB2A86AD429B08274824C98889D260D9159026741989D19",
            INIT_RAM_1F => X"48C0D04527CDF2031478C3CA2A02418F0A178864D51CA334C2434A633AA08A80",
            INIT_RAM_20 => X"04040404013403085049052444D1341C22016449404A14120D0117C8105851F2",
            INIT_RAM_21 => X"0CA0995511A0911A04200C5E11A440127043404C85412EA06194CACA80D04020",
            INIT_RAM_22 => X"75871C4508A52D19C51169487A4B5025A580117004820D85CD0401214D08602B",
            INIT_RAM_23 => X"419161A5DA0808D8488952531405314C104AA855594C1554115054A583370184",
            INIT_RAM_24 => X"0B04A1060A3268028A490414128C0935C115A1121861A5D1D9919219C602AA15",
            INIT_RAM_25 => X"140014B4027542430862A15431323005250502C85C9A028DD003542086012101",
            INIT_RAM_26 => X"22920D2480D24F3373742482BCE348523778D93C1202A154028C900829027C10",
            INIT_RAM_27 => X"01E34C2403B2B40308D1340842AD539B28384CE08E0A524020F0500E038ACC38",
            INIT_RAM_28 => X"0C080120DEE6F324070C11D1D190089034540B8C20BB0142C301430253244851",
            INIT_RAM_29 => X"15959D9D5D044404539AB9AA1801CC5516649DD35774C8C0006194C54002C01D",
            INIT_RAM_2A => X"86850600522132130A8A1A2A3A197577767657547446EA682015DC101AB99505",
            INIT_RAM_2B => X"76546C0911580045E104441A114045113460C8E0900317108BA29201082EA666",
            INIT_RAM_2C => X"44C11004013341D50474475455257214886EA6515959D9D30194CC2C5A268DA1",
            INIT_RAM_2D => X"026A01423448C808484056C2B0441E02493C2285F000C2008A240BC40404D104",
            INIT_RAM_2E => X"45917721B80E0020841514454953572144DD9955A0B016AAA060054565676408",
            INIT_RAM_2F => X"001D88D00D080152D1B54A457816361416214C6C11929D6E064B648744511574",
            INIT_RAM_30 => X"18036540DD1184050481121855611087214A52764012070D810DD5D3274851D8",
            INIT_RAM_31 => X"10A0A20B04546A311A448511722845063000EC0D0D8581C001627004D0605CC8",
            INIT_RAM_32 => X"064C21204D58014318C02A5E1711403C0F405134094A41305254C211DF0F0218",
            INIT_RAM_33 => X"59B676134820D0623498C889649B605341610802920A888C1362304D19713520",
            INIT_RAM_34 => X"3411166767243A45555941086D12404362221D920D2608DD8840367424840169",
            INIT_RAM_35 => X"02B3C32E107460623C700540D30CC0048CDC008CCDCF227C42F0033060010511",
            INIT_RAM_36 => X"7CC9700707078C924047089B005D4B043485314D220C11E378C157224059098B",
            INIT_RAM_37 => X"E01F0001C00841151116D5E0305CC1CBC010B89084018040C9104C97327A0216",
            INIT_RAM_38 => X"9FE803F7F510A0040D11F007402F3478E006CC0001B377504840440100448F28",
            INIT_RAM_39 => X"9BC04130626128E01EBD2261585582FD80B30100714E016841C506CC07DD583D",
            INIT_RAM_3A => X"05005003983225880911D1257660B45211D10D8195D1141C5C9454185458B8C8",
            INIT_RAM_3B => X"B216A194086821D07427705527C0000E60C89858585030F080C5591566A18216",
            INIT_RAM_3C => X"01C196419C6D526245CB093618906C921647F6709C48581310434C8562665140",
            INIT_RAM_3D => X"FFFFFFFFFFFFFFFFFFFFF26F0BFB518F50364F9AC9824B798DD8861F995A3460",
            INIT_RAM_3E => X"FFFFC09C931F19CB1F03C008D8D0035455C4D4C99C48140DCDDCD10E2390C562",
            INIT_RAM_3F => X"CCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"A8F9F2B492692201030004FC98B498CC2697475587CDD5746467675778D97857",
            INIT_RAM_01 => X"6603760570712DF1E06C55413D87DFCD34C541353446D375744E54E116735DE6",
            INIT_RAM_02 => X"3D63501F7174C716D661574803144DE534C783097DC00C44101ED3F373EE147F",
            INIT_RAM_03 => X"11614565051942A9586561D3088A903540E4350E24083AA8842CBBB0E03045C4",
            INIT_RAM_04 => X"100025902990190A07A079205C005106A8B682221A8805204C1850A025544891",
            INIT_RAM_05 => X"05D5D591155C10946200840658299A9DED199A29591918044344417112710C51",
            INIT_RAM_06 => X"86E144C28EC20ACE461020A22A20442210086A0243C002119952283ADD91D316",
            INIT_RAM_07 => X"4292A438EA9DC201A821A86D090E42864E0182D82114125E5A3BAAAAAAAB8AD2",
            INIT_RAM_08 => X"155534A64A6288B0922A28C88620881AC89909904820101A02B4423ACD01D468",
            INIT_RAM_09 => X"005062A2818081011E411AC40C46C0104219105E91E981D2B0F8F96181DDDD91",
            INIT_RAM_0A => X"5A625869C02AABA401C124A1069206A2C5BA418EC1D2662A20887850A8E52816",
            INIT_RAM_0B => X"1370C5011A42508200CF290036514588A5A6C72031080710AB114EDDE182493A",
            INIT_RAM_0C => X"FCD92280095995193C371072C1402AA66576714720E01D824A63E0A0AB39F02B",
            INIT_RAM_0D => X"586996B33F348E805EC14A44A7149949146A0650413700BA5A6194025D85C1BC",
            INIT_RAM_0E => X"6790440B390313934293A01F7C0084136424A02408293603667742438140469C",
            INIT_RAM_0F => X"C99DD03027DD49DC8DDC1C910701B092A4B64A95F1B304064444444446185284",
            INIT_RAM_10 => X"4AD8A828DAA2A8DE010492880376C0020CD922B393A39200A04C9324C0337438",
            INIT_RAM_11 => X"DD813AAB8B600DD82A17B28EC0EA808A0880273229248DA3A4A3242ECEA38107",
            INIT_RAM_12 => X"4D314689007005111115195F044687479246E01A07B8A24A9209451D9920B395",
            INIT_RAM_13 => X"C0446BC0420D82D0A0240A72F930051111151AC3900628AD8108809476E9A429",
            INIT_RAM_14 => X"3D4F42E9C06109512E7006AAAAA8040257C0042D043C4D4CB53D806727824005",
            INIT_RAM_15 => X"830D468C98CC9099288092A024A400AA405404F8C0036692830380AE9353C439",
            INIT_RAM_16 => X"61A990182C0EDB6DB5CA1846871CE39A21A2A1064981501ADC0926929106A187",
            INIT_RAM_17 => X"3C003BAEA483B0E0C3B7EDBB7888021C080947090A193934AC0CD23645659658",
            INIT_RAM_18 => X"6DDDDE1CDDD9DDE343C9C01F87EAA3BAA02ADB6A49248000CA9F03777C8E90F0",
            INIT_RAM_19 => X"04034A47F806A00CCC4CB052AC1ED428DA55315777489D2DE7009579424DF677",
            INIT_RAM_1A => X"86A90B2069A08962043536643644BB0A194C8ADE864D20CA344334330D001D00",
            INIT_RAM_1B => X"A0B70603000558265AD156092A628A288A16810DD954C5581A551D99DD03293A",
            INIT_RAM_1C => X"F8C1262A68921506808D4199DDDB6B3438083D0F60E0EA586F219682DB674732",
            INIT_RAM_1D => X"2561249921D30205A5C5CD199C22A22A2A8D288AB6168194988CE3B484DE1340",
            INIT_RAM_1E => X"24962581165595664A6298D9D1ADB08A663FB48A4C8DB6A992D8A36261809D95",
            INIT_RAM_1F => X"8F421965964AB24F04A0E3C3D029C2D5C3774046D188203409C9696A2672AA80",
            INIT_RAM_20 => X"32B2B2B20586CC00DB682595721C865716291729430036DA4A2DB7C9F7741293",
            INIT_RAM_21 => X"6DD01D1D1D3F1014C990289982666D808352722CDD99D9037748DDDD00EA9024",
            INIT_RAM_22 => X"4954044D4D11D91643114442A647740455421222070A51118D4018046E845A97",
            INIT_RAM_23 => X"6111DD11990944981C410A0A020080C05451101168249542550A00113C350554",
            INIT_RAM_24 => X"0BC0326403374C00F84CA0269A492DB4FC956C5844551152959C1A614D004404",
            INIT_RAM_25 => X"B0220A840149617141184046A07042A0A0A008C11DD905011A8802A211A8A8A8",
            INIT_RAM_26 => X"0C420DB6AA186B33437A302A800244A0378BEC800C084046A8CDD22AAC4B000E",
            INIT_RAM_27 => X"C10E43201466402A0002801605111846654570103D0DD2033F0E00810B404DC4",
            INIT_RAM_28 => X"15D04DB210197C10C713D951E14138A21640244000140002037800C04776442D",
            INIT_RAM_29 => X"5DD5DD5D91074A2AA7677777368180D10B442D10A47A000CC950664A904C102E",
            INIT_RAM_2A => X"0109AA328444446450F8343536267A77B77B77B47849DDD4DCD2ECD9377649FD",
            INIT_RAM_2B => X"555494C413A4904A81198427119042D2BB7F007200005050A01060002CA11111",
            INIT_RAM_2C => X"5B0D24EC4DB04D109496454250940044CA95555555555558229F04D8D5354D52",
            INIT_RAM_2D => X"8555C8B2168AD54D58D52C8D5376272104DC904A70044D42400A09C6D7A4E106",
            INIT_RAM_2E => X"60D834045C95404E09D0B4842D0B40045BD5D5D53D13A6AA909B975575575644",
            INIT_RAM_2F => X"D4104A005105719DD2BB634B5C083A18D7C1C498D2621947098A4505490D8378",
            INIT_RAM_30 => X"600B77579DDA884664CAD054DDD2181712B2407A81AA357E018D09EA3420D208",
            INIT_RAM_31 => X"2A424268C018941225C8099A4266398B270C944A828EC64301B3A0C4A414EC8A",
            INIT_RAM_32 => X"0AF0D2A44EE01209E0720DD59B0385516C2B92802A6A6C25A2A53D91572728E4",
            INIT_RAM_33 => X"DDBB762B4024E8923AE900A64A2B92A1A90910C973250C0722831C8E9A720A00",
            INIT_RAM_34 => X"3A0620A0AA2AB20982EA628C9A83A0A3A4022E964EB924EEA95ABAB920044B6E",
            INIT_RAM_35 => X"C7AC705A80785362AC70390A4260703A4C5703170107229C01F42F10B0000822",
            INIT_RAM_36 => X"1C997C1AC71909918A4A88281C914877452280A99140AD405402972380100DC0",
            INIT_RAM_37 => X"5C2710CE7C118D29D12DDDD4209C8E49C0689C4A961042909981A99726642A46",
            INIT_RAM_38 => X"667503B8B8EE7C3B8112701AC0C904908F2A0090C680786050C858C6724A4714",
            INIT_RAM_39 => X"21C0A2B0A2A3501002B2F037BCBFFC25A88C263390A8339C4242B60086E0D645",
            INIT_RAM_3A => X"082423146893196201E125B75468A73C1ADAD9CE9111E99C655CA5511C6A724C",
            INIT_RAM_3B => X"32664262099001DBBB3B7085050C8C51A24C2115511CC2400C80090008404044",
            INIT_RAM_3C => X"964CEC51A08F72F7394D108820D587B34F1CCF81C43110641561A4C282569960",
            INIT_RAM_3D => X"FFFFFFFFFFFFFFFFFFFFF2FC1730B20581988CB305030F8142000523BB510580",
            INIT_RAM_3E => X"FFFFC0BD04363043321F322024E08B3422CCCE422CE1F7C246E8E12E1360CDAC",
            INIT_RAM_3F => X"CCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1EE497BCFFCFBFFCFCFCCDCCFFCFFE8A0EDCABB9AD9FFEA9A8989A8AA8B9BB9A",
            INIT_RAM_01 => X"061406050401410105010044010410114115114045101441001015010504008A",
            INIT_RAM_02 => X"410E04504001102024064090101950004404141400155111541007F401AA4540",
            INIT_RAM_03 => X"C60E3AB838EEADAAAB2AB0C9A5990C161050340C5A403AAC0100000208452105",
            INIT_RAM_04 => X"982A68C8C2BA8A69AB9AB9AA828C0442AFA6EFB4B122406429EF3F8B4889BD26",
            INIT_RAM_05 => X"18E868E0022B6D3BB4DF7079C8EEAEACEECCE6CACACECB21B92ABACA843BCE00",
            INIT_RAM_06 => X"62A53270BC98B0707088AA9849973342ED2B937C2B07C9CCEEBB490C6CC2E8A0",
            INIT_RAM_07 => X"040FBF0C12E490F8FF8380042C9C1C961CFA784F83822A8CA043AAAAAAABE916",
            INIT_RAM_08 => X"022AB0BB0BB4D8B65ECAC319184359607B882EE818513D8F6318B60474B3496E",
            INIT_RAM_09 => X"CD852CACAAA3B8244E146A1B8E5830AEBA60C60EE0EE680278C8CA2A60CCCEE0",
            INIT_RAM_0A => X"20822096298A9881AAA82D9BE33F630CE4BB7A7C5B3622CAE5B2328626E6AD92",
            INIT_RAM_0B => X"E0B8E210240C032D3281F0CC800C8AA0861A2FAA38602FB9A4CCA68ACEAAAB98",
            INIT_RAM_0C => X"B200CADEA0022002804996CA060A9A8008800C8B53CA400F8BB308C8E0D2832E",
            INIT_RAM_0D => X"082082A080A2306A4ED80A80A96EEE3848B4D0A6BA0A820820820A62A2EB06C9",
            INIT_RAM_0E => X"92BD10AAE2E3A086140C0EACA0C2F986AEA300AEDB82D2CD1199090AE8840962",
            INIT_RAM_0F => X"ECC66DACA0AA3CA11CA10B0542CB81AAAE1AEA44BAC3985199911B91B8E19D31",
            INIT_RAM_10 => X"AA0D26232098A60265219AEA8409B2EBA76BBF0E2D2D1FC2BA5715C572D910AB",
            INIT_RAM_11 => X"223ABAABA8AA102181EBAA82AD026FF22BAEA83B49A31205298D852CF2ECA850",
            INIT_RAM_12 => X"963802E9AE8420066442244B912198A49A6B156B92A2BAEEB86220022BAAA000",
            INIT_RAM_13 => X"0E99AC528A300C032CC2588A0BAC200664422B0E0C2EBEA22EBA048891A4E384",
            INIT_RAM_14 => X"0C0370FFA2EBA66C0FF8B2AA2A9B23A912E321014581201C00402153ACA6372A",
            INIT_RAM_15 => X"B016D2F9690E4944081C16B090A6988088004A06F8CDB9BAE3B602622000C070",
            INIT_RAM_16 => X"2824A8E2EE38A28A2BA1CBB2ABE820688ACAD4E95460012845795AB8AAE9AE33",
            INIT_RAM_17 => X"3044AAAAAEBA418D052CCAB2AED658E3A0488862E1E3E2EEF0CE42AB332CB2CB",
            INIT_RAM_18 => X"A464ABB244A44AB90AEA0A85E17AAA00AE80A2AAABAEBA48E83C8DA22E929A02",
            INIT_RAM_19 => X"AD0A2AEC38EA223EB9F14F842ECEA123AECCEBBA223A44292E8BB3B39EAB1192",
            INIT_RAM_1A => X"AAD841692A4B91865AF07A20BBA0A01A8D0E804E18FBB4E86E1390A03B824408",
            INIT_RAM_1B => X"8528FAA38068806A8869101A26A492490A58962CC2AA288049882E88EE0A8840",
            INIT_RAM_1C => X"02996ACA9B1E5850B2FE1088EE492A91E0201A0680C0FA492A86184861B8DEAA",
            INIT_RAM_1D => X"723643EE20C99C1A287A54ECCBA4242A261622901A5896C2C8A69A499269B59A",
            INIT_RAM_1E => X"A1B2CCBC9A4A52BA7B1EC14CAE6A2E373882C1901198A28CC24B15A68292AEEB",
            INIT_RAM_1F => X"B88820861AEAAAABA0AE8AE81A62B22D1A21088AE2FEE8DA987B9B847B2E9808",
            INIT_RAM_20 => X"94949496208280C2492A86181C07082E9B41D1C92DE8924AAA861AEA112280B9",
            INIT_RAM_21 => X"08821A1A1A8187AB2EED91EC87B3984E350D0FCE88CC44AA223244AA72EAE8AA",
            INIT_RAM_22 => X"0A23F23C1ECCEE82FC8E330AA20B9080089682FBE8AA00001C1500C8BC228AA1",
            INIT_RAM_23 => X"9A8A44EE885A15872510F2F2FCDF3F2381AEE1CE23C5A2BC8AF0F2CCC0704AAA",
            INIT_RAM_24 => X"283AEBBB6E99BEDA061B7CB2CAA98A2BC52AA5A2A6882282A8A7882AF68BB873",
            INIT_RAM_25 => X"A4AD883A8A0A06062CC88409048416AF2F0F236CCAAAA21026D47C0ECCAF2F0F",
            INIT_RAM_26 => X"2AAC2492AA8A2AAEB633DC903AEAE380A3B0C77AE3678739ABA66D8067157AE2",
            INIT_RAM_27 => X"7EE2EFAA803BB4AF82D23CB210ECE43B308B81C80ADABAA3ACC2F23CA90BA832",
            INIT_RAM_28 => X"CE85BACEEE8EC072DEB8ACCCCECB8E2BD91C93E30893E948FA09CBE912ABA74A",
            INIT_RAM_29 => X"EA8EA8EACAB20A50B23A2A2B694BA3830E0C3830F2B3E3EA1EC87A3CC21A822C",
            INIT_RAM_2A => X"117E8AEC8784C4F0FA02A868687B33A32A32A32B33AEAAAFA182C3AF6AAB0B48",
            INIT_RAM_2B => X"B330BA3CBAB2BAEAEB9B2E6FBABAEA823AAC13F9F0033330B3B2500099233333",
            INIT_RAM_2C => X"B81825971A5FAACF303B333CCF33CB3251EEEECEECEECEE560341F36ADAB6ADB",
            INIT_RAM_2D => X"BEEC38A6F6188E18E18E2EFAEA2B2EAF2C3EC2EAD822BAFB0BC97B6D38A3CEB3",
            INIT_RAM_2E => X"8DA368B33A6632AAAC8F2033C8F23CB3308E8E8E81BCB00014BC72BB2BB2BA97",
            INIT_RAM_2F => X"A3CF38F2CCB30CC882B28A0A3E88FAE3AD372DCFAB34DB2EACD27CB3ACDA36B3",
            INIT_RAM_30 => X"48AA22304A86833B3A74AB328882EACE8728FB3A1E6CEB0C1EBAFCE063C580F5",
            INIT_RAM_31 => X"EEDA868E23ED8D8F6BA178AE86AB4AC8694EA13838383853B42E14E183C181D2",
            INIT_RAM_32 => X"8BC1AE330DA1EA2B3ADB68822DA88B7B707C8ECC9290D1EA842B8ACCECAD8D32",
            INIT_RAM_33 => X"A8CEA37688B0D38C34AE53220B2B8C0C9A2EB25AEA63613EBB95FAEE8EEB88CC",
            INIT_RAM_34 => X"34C120407BCAE80481AAB21BAA0E3F03FB522C1B0D2860DE8E4028B04B393A33",
            INIT_RAM_35 => X"C5E2C6CECB338E84B2E89BE1D991E89B61EE89B81EBFB8B603F81F62F0088812",
            INIT_RAM_36 => X"F6CCE0ABEEABACCBAB0BEEEEB2CAD366FC82FC96DB210AEA3E16EEBA801F1FC2",
            INIT_RAM_37 => X"EEEDBAEAE09B282CAC288AAEBBBAEAB3E267BE3ACDA70ABACC049EEEBB3853B3",
            INIT_RAM_38 => X"9350034040E0F09BAAC2F8ABA26FA0BAE3BBA1BAEEEA328FB213B2EECB0B6DBE",
            INIT_RAM_39 => X"2409BEEE0F2A212006BF337A7771B63CF2E06CBA842EBBBEE6102BA1390261E2",
            INIT_RAM_3A => X"8A6303802EBBAA2AA4A82800230D37B64E0200AE0800200AE00AE0000E243AEE",
            INIT_RAM_3B => X"9BBB87B52CC22424B3C8151A5AE78E00BAEEE00006680EB821B5515559858910",
            INIT_RAM_3C => X"106001104650002000698401920514004819081904200AEA802BAEE2DB8AECAA",
            INIT_RAM_3D => X"FFFFFFFFFFFFFFFFFFFFF0209044092FF901500EE46EE0146042FF8400049148",
            INIT_RAM_3E => X"FFFFE80FEF95AEEE91AA09B101FA6F6102DAD2D02D8B3050346DFB4E8F72D19E",
            INIT_RAM_3F => X"CCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_2_AD_i
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 2,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"DF75D79F7DD75CCCFEEEECEDFFCEEEFE0FDFDDEDCCFDDCDDCDFECCEEEDFCFCDC",
            INIT_RAM_01 => X"565776575D57575755D5D7575757577575D55D57555DD7575D5D755D5D5D75E7",
            INIT_RAM_02 => X"555055555555552565565595D7595D7575D75D75D75D75D75D75D6ADD7AAD5D7",
            INIT_RAM_03 => X"8ACA9E8B2A728EEBA9AE8A6C1F848C3A30E82A08E8EC2FF85540050050554555",
            INIT_RAM_04 => X"D00EA5D0FAE3AB8F36F36F34524ACCAD9CE9EC33A624ACCAD2798847FBBAAFAA",
            INIT_RAM_05 => X"2A6A5A6AAAA32FDDFF661C947CA7A2B6D66652EA6A666A26C1B8D3DE0ABBC8EE",
            INIT_RAM_06 => X"C23227F7E7E3F33333E0B4F03F3999B166296FDB2D4D886666D32A0A666A6F2B",
            INIT_RAM_07 => X"8DCCC3082FA43BFECF32FFA62A23233A331473633262E56D64CD3FFFFFFF0D7F",
            INIT_RAM_08 => X"AAAE1859859B68BD3AAAA32B88E32B2F3AAA2667882C2BEB3ADFBF0BF7F26B71",
            INIT_RAM_09 => X"8CCCEBABD307A6222E3025BD08BB3330D3ECC9ED6ED616A2B8E4E59B0A66666A",
            INIT_RAM_0A => X"A691E7630C096863E386AFF23AF33ACFEA9CC4FFCD6EAABAA3ADB58CFC4A2D28",
            INIT_RAM_0B => X"FDF08F2EDABBAEDCE2C4CCF8AA8FBB069A6B4E3820ECCC3AB566EAA84AE38F29",
            INIT_RAM_0C => X"D52C8FFE1AAAAEEAD4E88F5D498BA96AAAAA8FB8C2D1AA898D825C9CA38F92B1",
            INIT_RAM_0D => X"E79A6971D4823BB8AEF78EB8E8B0662CBB488EB0D3DE0C69A69E7B02E74D4F5F",
            INIT_RAM_0E => X"98F88897CF42314EEECEDE3DE48CBC0EBCA3B338FF3FDFF99999898827CBB4B0",
            INIT_RAM_0F => X"4AAAAE28B1AA27A327A2BA8CAE8B53E0785BCAAAF3520C89480085885040B8D8",
            INIT_RAM_10 => X"992FFC2326F0BC22222FF38D08C4A2E34C4E1CDCDEDEDCCCE1AAEABAA2F2A8AB",
            INIT_RAM_11 => X"AA3673FF04F43322341082F74F3FC6BF2B8E3123FF23238ED73E131DE339D08C",
            INIT_RAM_12 => X"0423BB0F110CCEEAA22EEAAF2A9AAAB5F3CC432C08BCE3C2E0CD5EEAAE38B1AA",
            INIT_RAM_13 => X"4DAAB5FBC2EAFBAEDFB23BC35F0CCEE22AAEEF4CCCCD34E7CF38C87B98262336",
            INIT_RAM_14 => X"0A8230CBC2D34AAA0AC09BFFBFE723E2ABC32301551545500555455479E23A2C",
            INIT_RAM_15 => X"75356163AF48A6B910C8CAC328B8C0990BFCFB52E48100E3023CCCA1BDE0B82A",
            INIT_RAM_16 => X"965AE0DCDE15A69A6B8665D9B6AC7DAD1D9DB9B7FA2FF3E2577829C1E1B7651B",
            INIT_RAM_17 => X"24FC8820B8F312BC4EF9DAB6BC323BF78C87B8CFEDEFCDB4D488626AA69A69A6",
            INIT_RAM_18 => X"A545AF3865A65AF188EE48AFABE9F3569E19A6A78F38F0AC89314DAABCC54B52",
            INIT_RAM_19 => X"9F330BCF78D0B22EFBA2028FFEAEA223B2AAE2AAAAB8B62F6F0AAA128B8E5516",
            INIT_RAM_1A => X"5B1C9FFE1A27BE8EE8DCDEA89998B1334288A26E33ED3888B42218B12D0CA630",
            INIT_RAM_1B => X"8AE82B82029AACAA4466AB2A12ABAEBACAABAA266EABCAAC84AAA6AA6607A8CD",
            INIT_RAM_1C => X"520BA6BA4ACEE8EFA2373BAA66659F1BCCCC2A0A9090A9A69F1A698965B17F3B",
            INIT_RAM_1D => X"EEFEA3AB2A6C1F29AA69F76AAD2AEB16111422AFDAABAAA2A8B0F31FB26F3D8B",
            INIT_RAM_1E => X"A89AA6A66AA9AA6AE2388F7A96A9B4322BD752BB32BA6A7AA26ADDAAFAA2B62F",
            INIT_RAM_1F => X"B5C1E79A6BCAF38F1ABCF3CD4AFAF22F6AA98AEA7A30E0D9FBA96960A22A2888",
            INIT_RAM_20 => X"6B6B6B692E79C4CCA69E1A6BABEA79ED2B26AABAAE88A9A78F1A6BCE6AB068F2",
            INIT_RAM_21 => X"AAA22A2A2AD48DDB8AAE23AACAAA6A0CFDCDCEBEAAAA6626AAB0AAAA32E5D0B8",
            INIT_RAM_22 => X"8AABFC37376666A2FF0DD989AAA9A8AAAABD6AC21896AAAA2732B8AA4D556FD9",
            INIT_RAM_23 => X"4AAAAA66AA2B32B2B32B6E6CDB06FFCFB3B6726511BC2A5BA96C6266C4DCEEAA",
            INIT_RAM_24 => X"2F7CE2AB8E2AB4E3522928A9A78E1A6B1AEAEAAEBCAAAAA1AA9AA90AFA499C99",
            INIT_RAM_25 => X"689E09B8498D8DCDD666CAA44ECECC66E6D623C66AAE1B2A91FA9A4E666AEADA",
            INIT_RAM_26 => X"26CE2A6995A69F2AAAF6AC86F4E3C3332BB1DB34F789C994678AAE19AA2AF4F5",
            INIT_RAM_27 => X"8AE7CF387BAA989D0C62589B2E66539AABBBD3E0DAFAF38235E6623E198B8F78",
            INIT_RAM_28 => X"AAA23B3EAAAAE4F42D35AA9ADAD35EA7E248ABC330ABC48AF3D88BC48AAB0ABA",
            INIT_RAM_29 => X"9AA9AA9AA96A8BCC6AAAAAA8E88B02A30A8C2A30AA74A3BA48E06ACFA23AA21D",
            INIT_RAM_2A => X"202A8FF04A8888A89B526CECECEEB6AB6AB6AB6AB6999993B2A1DEB32222071A",
            INIT_RAM_2B => X"9998B47D3AB074EAD3AB4EAE3AB4EAAA5EB503E0482B0B098B1948024FD11113",
            INIT_RAM_2C => X"BD3A9000290E9AA6AA2AA69AA6A98999F695556966966960A8753C70AC2B0AC2",
            INIT_RAM_2D => X"E8882080DB20BA3BA3BA2EBBD2AC2E1F4F70A2EAE009FBD28B843B8D7D50DA6A",
            INIT_RAM_2E => X"A6A9A899B8AA32A29AA6AA29AA6A9899BDA6A6A6D4B128003DBDAAEAAEAAEACC",
            INIT_RAM_2F => X"BC96FB626667DAAAA236AA8AB848B8A3AC7F4E8FA6BFAA2E1AFEA8AA9A6A9A12",
            INIT_RAM_30 => X"889AAABD6AAA26AAB02BA6B8A898A9AD03EAC2BA08B1EBDD2A3B6B6CEDB3B863",
            INIT_RAM_31 => X"31E2C21F50AFBE0FEF803AB2B627DB08218893333B333B220DCCD88333A332CE",
            INIT_RAM_32 => X"CB53A2EA8E20822E74F0AAAAAD3A81B1B5B9A3348240D42188EB5AA9AF1E1E70",
            INIT_RAM_33 => X"AAE6AB92A8A8EC8E3B2A03AA8C2B48C04A2C34FBE3EF803F3880FCE2AEF3988E",
            INIT_RAM_34 => X"38C220A0878F0A09822AC203A2CCFCE3AACE8DAA8EC8ECE4BAAFC474AC0C2EB9",
            INIT_RAM_35 => X"4860694226B68E8970F0AB86E1A3F0AB40AD0ABD3A7C3AB803F40F0170248822",
            INIT_RAM_36 => X"B4AAF4AB4F2B4AA7468B4EEF34AACEAAA8933E46D382BAE2B825AF3B8084BD65",
            INIT_RAM_37 => X"AE6E34E6D4BBCAAAAA2AAAAD3ABCEAFB02E0B861527ECAB4AAC84AAF2AACEEAA",
            INIT_RAM_38 => X"2BC801C6C6C5E4AB46A2C0ABC2AF18B4D79BC074E6F1B582B406B4E6D28B4E38",
            INIT_RAM_39 => X"6767C33CC8F6F3F0269651935297169311F41D398ADD3AB8EA2B6BC06B1B6909",
            INIT_RAM_3A => X"88EB723BB0E3999B422A26489AAFEBE2222622E62A22622EA22EE2222E2ABB8E",
            INIT_RAM_3B => X"C199CDDA26622210F78CB8CBCB4388EEC38E6AAAA22C4ED0C3F320CCA8CCC888",
            INIT_RAM_3C => X"554555515455500555411555145554015151515154122E6D08BAB8EAD1EA72B4",
            INIT_RAM_3D => X"FFFFFFFFFFFFFFFFFFFFF0051555514001555500054005554554001500551550",
            INIT_RAM_3E => X"FFFFD401551515451515444332C113E330F9F9F30F9D71F737CEC3FC0F62FAAE",
            INIT_RAM_3F => X"CCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_3_AD_i
        );

end Behavioral; --basicRom
