//Copyright (C)2014-2021 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8
//Part Number: GW1NSR-LV4CQN48PC7/I6
//Device: GW1NSR-4C
//Created Time: Sun Sep 12 19:16:18 2021

module basicRom (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hEA460278D7349FCC8FD0C210FCF5C8ED2D2C0B0820DDC1AEBE9B9F88C606BB59;
defparam prom_inst_0.INIT_RAM_01 = 256'h40CEB093694CD0BC987C919C705C1ACCD6A469FDB3699B3C41650494406B8913;
defparam prom_inst_0.INIT_RAM_02 = 256'hC4130ED7BE3EBA0140D82423F462393521927FC1F0A9FC6ADE49BC6B26E7133A;
defparam prom_inst_0.INIT_RAM_03 = 256'h4180544EC952702DD16640DB0084B19DC745DD6605155008D6A49F9090BA49B3;
defparam prom_inst_0.INIT_RAM_04 = 256'hF0C4927300312441151113002211522008042722D02214020849536226E19406;
defparam prom_inst_0.INIT_RAM_05 = 256'h4C0159D8585CD88A90D52B14230D92D1D1DDD2491D5D99402138F18E20B8000E;
defparam prom_inst_0.INIT_RAM_06 = 256'h4D0D0C414541C1C50DE080102122594195094314093150858530093440D0D710;
defparam prom_inst_0.INIT_RAM_07 = 256'h614240249085C18044110B840801010D0D0009181100E01D10376AAAAAAB4220;
defparam prom_inst_0.INIT_RAM_08 = 256'h5853046765545050324A4809150C0990C9E94A53641018060D1B902401011810;
defparam prom_inst_0.INIT_RAM_09 = 256'h210264A4024490495D89500F00010208F104201D9DD505118991518A80D850D8;
defparam prom_inst_0.INIT_RAM_0A = 256'hD04113438A0429645345141301120102CCB4000D08336A4A4090746244DC1632;
defparam prom_inst_0.INIT_RAM_0B = 256'h1870028DD074DD20D8012734036036414D07CE2402248F1078854D55D1920F14;
defparam prom_inst_0.INIT_RAM_0C = 256'h8068208E00D850DDA302B209308914214343403504D00D121540004148074C11;
defparam prom_inst_0.INIT_RAM_0D = 256'h13413400A282C194DD4047756608A5030B432474F1890804D04D068D80833080;
defparam prom_inst_0.INIT_RAM_0E = 256'h7772988207C0280390404E1C9308CD107C1412244C900434B7840388A0A37438;
defparam prom_inst_0.INIT_RAM_0F = 256'h841C902404C9CD9400C8593326630CB22437CD0D33402A17569A65555A694156;
defparam prom_inst_0.INIT_RAM_10 = 256'h48A8841062124495AC080080336490218CC923407370730820D9364D90B32406;
defparam prom_inst_0.INIT_RAM_11 = 256'h85C936AB8280CD9C100341100C5045880A820402202C4980485F005D09040206;
defparam prom_inst_0.INIT_RAM_12 = 256'h0C003983222080E86850D0D321A443BC00CB08D6247023CDD32480D0D321400D;
defparam prom_inst_0.INIT_RAM_13 = 256'h32A1544CF2D9345D134A88E1CD0080D85850D030708C0C634F001043441D9C9D;
defparam prom_inst_0.INIT_RAM_14 = 256'h6755C44B84C000D146F138008020205034CC0024931E8C6C91BB46070C81C508;
defparam prom_inst_0.INIT_RAM_15 = 256'h64CD0D00EA00D4DD597372423470A1480B8A3A8243330092801048AD98177511;
defparam prom_inst_0.INIT_RAM_16 = 256'h4D8483040C101149378091940A1020DE03405109CDCE28EAE0CB10F080090597;
defparam prom_inst_0.INIT_RAM_17 = 256'h0334041164E0CC523274D93754C0C5F081043727340427143300D10447491413;
defparam prom_inst_0.INIT_RAM_18 = 256'h4515D53C15DD595100C804DF6790D0820E0893628D24E01008BC13B24CD0128A;
defparam prom_inst_0.INIT_RAM_19 = 256'h80210B4F3636868EC55030B20C1D20501286A2161868ED112C03447772CD1756;
defparam prom_inst_0.INIT_RAM_1A = 256'h0535140499049042761422780B546CC1508086DDC185300B14403880C508DA20;
defparam prom_inst_0.INIT_RAM_1B = 256'h50450640000411325652144C9264924906449D085105C41124C90DC985012724;
defparam prom_inst_0.INIT_RAM_1C = 256'h820B364A49224634904C01DA96934F1204815D6645466013470D0400D2440C13;
defparam prom_inst_0.INIT_RAM_1D = 256'h39B0448E10DB20C18545064DAC26241250081E9016449DA2D06C630C9056326A;
defparam prom_inst_0.INIT_RAM_1E = 256'h84764994149514648AB2A86AD429B08274824C98889D260D9159026741989D19;
defparam prom_inst_0.INIT_RAM_1F = 256'h48C0D04527CDF2031478C3CA2A02418F0A178864D51CA334C2434A633AA08A80;
defparam prom_inst_0.INIT_RAM_20 = 256'h04040404013403085049052444D1341C22016449404A14120D0117C8105851F2;
defparam prom_inst_0.INIT_RAM_21 = 256'h0CA0995511A0911A04200C5E11A440127043404C85412EA06194CACA80D04020;
defparam prom_inst_0.INIT_RAM_22 = 256'h75871C4508A52D19C51169487A4B5025A580117004820D85CD0401214D08602B;
defparam prom_inst_0.INIT_RAM_23 = 256'h419161A5DA0808D8488952531405314C104AA855594C1554115054A583370184;
defparam prom_inst_0.INIT_RAM_24 = 256'h0B04A1060A3268028A490414128C0935C115A1121861A5D1D9919219C602AA15;
defparam prom_inst_0.INIT_RAM_25 = 256'h140014B4027542430862A15431323005250502C85C9A028DD003542086012101;
defparam prom_inst_0.INIT_RAM_26 = 256'h22920D2480D24F3373742482BCE348523778D93C1202A154028C900829027C10;
defparam prom_inst_0.INIT_RAM_27 = 256'h01E34C2403B2B40308D1340842AD539B28384CE08E0A524020F0500E038ACC38;
defparam prom_inst_0.INIT_RAM_28 = 256'h0C080120DEE6F324070C11D1D190089034540B8C20BB0142C301430253244851;
defparam prom_inst_0.INIT_RAM_29 = 256'h15959D9D5D044404539AB9AA1801CC5516649DD35774C8C0006194C54002C01D;
defparam prom_inst_0.INIT_RAM_2A = 256'h86850600522132130A8A1A2A3A197577767657547446EA682015DC101AB99505;
defparam prom_inst_0.INIT_RAM_2B = 256'h76546C0911580045E104441A114045113460C8E0900317108BA29201082EA666;
defparam prom_inst_0.INIT_RAM_2C = 256'h44C11004013341D50474475455257214886EA6515959D9D30194CC2C5A268DA1;
defparam prom_inst_0.INIT_RAM_2D = 256'h026A01423448C808484056C2B0441E02493C2285F000C2008A240BC40404D104;
defparam prom_inst_0.INIT_RAM_2E = 256'h45917721B80E0020841514454953572144DD9955A0B016AAA060054565676408;
defparam prom_inst_0.INIT_RAM_2F = 256'h001D88D00D080152D1B54A457816361416214C6C11929D6E064B648744511574;
defparam prom_inst_0.INIT_RAM_30 = 256'h18036540DD1184050481121855611087214A52764012070D810DD5D3274851D8;
defparam prom_inst_0.INIT_RAM_31 = 256'h10A0A20B04546A311A448511722845063000EC0D0D8581C001627004D0605CC8;
defparam prom_inst_0.INIT_RAM_32 = 256'h064C21204D58014318C02A5E1711403C0F405134094A41305254C211DF0F0218;
defparam prom_inst_0.INIT_RAM_33 = 256'h59B676134820D0623498C889649B605341610802920A888C1362304D19713520;
defparam prom_inst_0.INIT_RAM_34 = 256'h3411166767243A45555941086D12404362221D920D2608DD8840367424840169;
defparam prom_inst_0.INIT_RAM_35 = 256'h02B3C32E107460623C700540D30CC0048CDC008CCDCF227C42F0033060010511;
defparam prom_inst_0.INIT_RAM_36 = 256'h7CC9700707078C924047089B005D4B043485314D220C11E378C157224059098B;
defparam prom_inst_0.INIT_RAM_37 = 256'hE01F0001C00841151116D5E0305CC1CBC010B89084018040C9104C97327A0216;
defparam prom_inst_0.INIT_RAM_38 = 256'h9FE803F7F510A0040D11F007402F3478E006CC0001B377504840440100448F28;
defparam prom_inst_0.INIT_RAM_39 = 256'h9BC04130626128E01EBD2261585582FD80B30100714E016841C506CC07DD583D;
defparam prom_inst_0.INIT_RAM_3A = 256'h05005003983225880911D1257660B45211D10D8195D1141C5C9454185458B8C8;
defparam prom_inst_0.INIT_RAM_3B = 256'hB216A194086821D07427705527C0000E60C89858585030F080C5591566A18216;
defparam prom_inst_0.INIT_RAM_3C = 256'h01C196419C6D526245CB093618906C921647F6709C48581310434C8562665140;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFF26F0BFB518F50364F9AC9824B798DD8861F995A3460;
defparam prom_inst_0.INIT_RAM_3E = 256'hFFFFC09C931F19CB1F03C008D8D0035455C4D4C99C48140DCDDCD10E2390C562;
defparam prom_inst_0.INIT_RAM_3F = 256'hCCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hA8F9F2B492692201030004FC98B498CC2697475587CDD5746467675778D97857;
defparam prom_inst_1.INIT_RAM_01 = 256'h6603760570712DF1E06C55413D87DFCD34C541353446D375744E54E116735DE6;
defparam prom_inst_1.INIT_RAM_02 = 256'h3D63501F7174C716D661574803144DE534C783097DC00C44101ED3F373EE147F;
defparam prom_inst_1.INIT_RAM_03 = 256'h11614565051942A9586561D3088A903540E4350E24083AA8842CBBB0E03045C4;
defparam prom_inst_1.INIT_RAM_04 = 256'h100025902990190A07A079205C005106A8B682221A8805204C1850A025544891;
defparam prom_inst_1.INIT_RAM_05 = 256'h05D5D591155C10946200840658299A9DED199A29591918044344417112710C51;
defparam prom_inst_1.INIT_RAM_06 = 256'h86E144C28EC20ACE461020A22A20442210086A0243C002119952283ADD91D316;
defparam prom_inst_1.INIT_RAM_07 = 256'h4292A438EA9DC201A821A86D090E42864E0182D82114125E5A3BAAAAAAAB8AD2;
defparam prom_inst_1.INIT_RAM_08 = 256'h155534A64A6288B0922A28C88620881AC89909904820101A02B4423ACD01D468;
defparam prom_inst_1.INIT_RAM_09 = 256'h005062A2818081011E411AC40C46C0104219105E91E981D2B0F8F96181DDDD91;
defparam prom_inst_1.INIT_RAM_0A = 256'h5A625869C02AABA401C124A1069206A2C5BA418EC1D2662A20887850A8E52816;
defparam prom_inst_1.INIT_RAM_0B = 256'h1370C5011A42508200CF290036514588A5A6C72031080710AB114EDDE182493A;
defparam prom_inst_1.INIT_RAM_0C = 256'hFCD92280095995193C371072C1402AA66576714720E01D824A63E0A0AB39F02B;
defparam prom_inst_1.INIT_RAM_0D = 256'h586996B33F348E805EC14A44A7149949146A0650413700BA5A6194025D85C1BC;
defparam prom_inst_1.INIT_RAM_0E = 256'h6790440B390313934293A01F7C0084136424A02408293603667742438140469C;
defparam prom_inst_1.INIT_RAM_0F = 256'hC99DD03027DD49DC8DDC1C910701B092A4B64A95F1B304064444444446185284;
defparam prom_inst_1.INIT_RAM_10 = 256'h4AD8A828DAA2A8DE010492880376C0020CD922B393A39200A04C9324C0337438;
defparam prom_inst_1.INIT_RAM_11 = 256'hDD813AAB8B600DD82A17B28EC0EA808A0880273229248DA3A4A3242ECEA38107;
defparam prom_inst_1.INIT_RAM_12 = 256'h4D314689007005111115195F044687479246E01A07B8A24A9209451D9920B395;
defparam prom_inst_1.INIT_RAM_13 = 256'hC0446BC0420D82D0A0240A72F930051111151AC3900628AD8108809476E9A429;
defparam prom_inst_1.INIT_RAM_14 = 256'h3D4F42E9C06109512E7006AAAAA8040257C0042D043C4D4CB53D806727824005;
defparam prom_inst_1.INIT_RAM_15 = 256'h830D468C98CC9099288092A024A400AA405404F8C0036692830380AE9353C439;
defparam prom_inst_1.INIT_RAM_16 = 256'h61A990182C0EDB6DB5CA1846871CE39A21A2A1064981501ADC0926929106A187;
defparam prom_inst_1.INIT_RAM_17 = 256'h3C003BAEA483B0E0C3B7EDBB7888021C080947090A193934AC0CD23645659658;
defparam prom_inst_1.INIT_RAM_18 = 256'h6DDDDE1CDDD9DDE343C9C01F87EAA3BAA02ADB6A49248000CA9F03777C8E90F0;
defparam prom_inst_1.INIT_RAM_19 = 256'h04034A47F806A00CCC4CB052AC1ED428DA55315777489D2DE7009579424DF677;
defparam prom_inst_1.INIT_RAM_1A = 256'h86A90B2069A08962043536643644BB0A194C8ADE864D20CA344334330D001D00;
defparam prom_inst_1.INIT_RAM_1B = 256'hA0B70603000558265AD156092A628A288A16810DD954C5581A551D99DD03293A;
defparam prom_inst_1.INIT_RAM_1C = 256'hF8C1262A68921506808D4199DDDB6B3438083D0F60E0EA586F219682DB674732;
defparam prom_inst_1.INIT_RAM_1D = 256'h2561249921D30205A5C5CD199C22A22A2A8D288AB6168194988CE3B484DE1340;
defparam prom_inst_1.INIT_RAM_1E = 256'h24962581165595664A6298D9D1ADB08A663FB48A4C8DB6A992D8A36261809D95;
defparam prom_inst_1.INIT_RAM_1F = 256'h8F421965964AB24F04A0E3C3D029C2D5C3774046D188203409C9696A2672AA80;
defparam prom_inst_1.INIT_RAM_20 = 256'h32B2B2B20586CC00DB682595721C865716291729430036DA4A2DB7C9F7741293;
defparam prom_inst_1.INIT_RAM_21 = 256'h6DD01D1D1D3F1014C990289982666D808352722CDD99D9037748DDDD00EA9024;
defparam prom_inst_1.INIT_RAM_22 = 256'h4954044D4D11D91643114442A647740455421222070A51118D4018046E845A97;
defparam prom_inst_1.INIT_RAM_23 = 256'h6111DD11990944981C410A0A020080C05451101168249542550A00113C350554;
defparam prom_inst_1.INIT_RAM_24 = 256'h0BC0326403374C00F84CA0269A492DB4FC956C5844551152959C1A614D004404;
defparam prom_inst_1.INIT_RAM_25 = 256'hB0220A840149617141184046A07042A0A0A008C11DD905011A8802A211A8A8A8;
defparam prom_inst_1.INIT_RAM_26 = 256'h0C420DB6AA186B33437A302A800244A0378BEC800C084046A8CDD22AAC4B000E;
defparam prom_inst_1.INIT_RAM_27 = 256'hC10E43201466402A0002801605111846654570103D0DD2033F0E00810B404DC4;
defparam prom_inst_1.INIT_RAM_28 = 256'h15D04DB210197C10C713D951E14138A21640244000140002037800C04776442D;
defparam prom_inst_1.INIT_RAM_29 = 256'h5DD5DD5D91074A2AA7677777368180D10B442D10A47A000CC950664A904C102E;
defparam prom_inst_1.INIT_RAM_2A = 256'h0109AA328444446450F8343536267A77B77B77B47849DDD4DCD2ECD9377649FD;
defparam prom_inst_1.INIT_RAM_2B = 256'h555494C413A4904A81198427119042D2BB7F007200005050A01060002CA11111;
defparam prom_inst_1.INIT_RAM_2C = 256'h5B0D24EC4DB04D109496454250940044CA95555555555558229F04D8D5354D52;
defparam prom_inst_1.INIT_RAM_2D = 256'h8555C8B2168AD54D58D52C8D5376272104DC904A70044D42400A09C6D7A4E106;
defparam prom_inst_1.INIT_RAM_2E = 256'h60D834045C95404E09D0B4842D0B40045BD5D5D53D13A6AA909B975575575644;
defparam prom_inst_1.INIT_RAM_2F = 256'hD4104A005105719DD2BB634B5C083A18D7C1C498D2621947098A4505490D8378;
defparam prom_inst_1.INIT_RAM_30 = 256'h600B77579DDA884664CAD054DDD2181712B2407A81AA357E018D09EA3420D208;
defparam prom_inst_1.INIT_RAM_31 = 256'h2A424268C018941225C8099A4266398B270C944A828EC64301B3A0C4A414EC8A;
defparam prom_inst_1.INIT_RAM_32 = 256'h0AF0D2A44EE01209E0720DD59B0385516C2B92802A6A6C25A2A53D91572728E4;
defparam prom_inst_1.INIT_RAM_33 = 256'hDDBB762B4024E8923AE900A64A2B92A1A90910C973250C0722831C8E9A720A00;
defparam prom_inst_1.INIT_RAM_34 = 256'h3A0620A0AA2AB20982EA628C9A83A0A3A4022E964EB924EEA95ABAB920044B6E;
defparam prom_inst_1.INIT_RAM_35 = 256'hC7AC705A80785362AC70390A4260703A4C5703170107229C01F42F10B0000822;
defparam prom_inst_1.INIT_RAM_36 = 256'h1C997C1AC71909918A4A88281C914877452280A99140AD405402972380100DC0;
defparam prom_inst_1.INIT_RAM_37 = 256'h5C2710CE7C118D29D12DDDD4209C8E49C0689C4A961042909981A99726642A46;
defparam prom_inst_1.INIT_RAM_38 = 256'h667503B8B8EE7C3B8112701AC0C904908F2A0090C680786050C858C6724A4714;
defparam prom_inst_1.INIT_RAM_39 = 256'h21C0A2B0A2A3501002B2F037BCBFFC25A88C263390A8339C4242B60086E0D645;
defparam prom_inst_1.INIT_RAM_3A = 256'h082423146893196201E125B75468A73C1ADAD9CE9111E99C655CA5511C6A724C;
defparam prom_inst_1.INIT_RAM_3B = 256'h32664262099001DBBB3B7085050C8C51A24C2115511CC2400C80090008404044;
defparam prom_inst_1.INIT_RAM_3C = 256'h964CEC51A08F72F7394D108820D587B34F1CCF81C43110641561A4C282569960;
defparam prom_inst_1.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFF2FC1730B20581988CB305030F8142000523BB510580;
defparam prom_inst_1.INIT_RAM_3E = 256'hFFFFC0BD04363043321F322024E08B3422CCCE422CE1F7C246E8E12E1360CDAC;
defparam prom_inst_1.INIT_RAM_3F = 256'hCCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h1EE497BCFFCFBFFCFCFCCDCCFFCFFE8A0EDCABB9AD9FFEA9A8989A8AA8B9BB9A;
defparam prom_inst_2.INIT_RAM_01 = 256'h061406050401410105010044010410114115114045101441001015010504008A;
defparam prom_inst_2.INIT_RAM_02 = 256'h410E04504001102024064090101950004404141400155111541007F401AA4540;
defparam prom_inst_2.INIT_RAM_03 = 256'hC60E3AB838EEADAAAB2AB0C9A5990C161050340C5A403AAC0100000208452105;
defparam prom_inst_2.INIT_RAM_04 = 256'h982A68C8C2BA8A69AB9AB9AA828C0442AFA6EFB4B122406429EF3F8B4889BD26;
defparam prom_inst_2.INIT_RAM_05 = 256'h18E868E0022B6D3BB4DF7079C8EEAEACEECCE6CACACECB21B92ABACA843BCE00;
defparam prom_inst_2.INIT_RAM_06 = 256'h62A53270BC98B0707088AA9849973342ED2B937C2B07C9CCEEBB490C6CC2E8A0;
defparam prom_inst_2.INIT_RAM_07 = 256'h040FBF0C12E490F8FF8380042C9C1C961CFA784F83822A8CA043AAAAAAABE916;
defparam prom_inst_2.INIT_RAM_08 = 256'h022AB0BB0BB4D8B65ECAC319184359607B882EE818513D8F6318B60474B3496E;
defparam prom_inst_2.INIT_RAM_09 = 256'hCD852CACAAA3B8244E146A1B8E5830AEBA60C60EE0EE680278C8CA2A60CCCEE0;
defparam prom_inst_2.INIT_RAM_0A = 256'h20822096298A9881AAA82D9BE33F630CE4BB7A7C5B3622CAE5B2328626E6AD92;
defparam prom_inst_2.INIT_RAM_0B = 256'hE0B8E210240C032D3281F0CC800C8AA0861A2FAA38602FB9A4CCA68ACEAAAB98;
defparam prom_inst_2.INIT_RAM_0C = 256'hB200CADEA0022002804996CA060A9A8008800C8B53CA400F8BB308C8E0D2832E;
defparam prom_inst_2.INIT_RAM_0D = 256'h082082A080A2306A4ED80A80A96EEE3848B4D0A6BA0A820820820A62A2EB06C9;
defparam prom_inst_2.INIT_RAM_0E = 256'h92BD10AAE2E3A086140C0EACA0C2F986AEA300AEDB82D2CD1199090AE8840962;
defparam prom_inst_2.INIT_RAM_0F = 256'hECC66DACA0AA3CA11CA10B0542CB81AAAE1AEA44BAC3985199911B91B8E19D31;
defparam prom_inst_2.INIT_RAM_10 = 256'hAA0D26232098A60265219AEA8409B2EBA76BBF0E2D2D1FC2BA5715C572D910AB;
defparam prom_inst_2.INIT_RAM_11 = 256'h223ABAABA8AA102181EBAA82AD026FF22BAEA83B49A31205298D852CF2ECA850;
defparam prom_inst_2.INIT_RAM_12 = 256'h963802E9AE8420066442244B912198A49A6B156B92A2BAEEB86220022BAAA000;
defparam prom_inst_2.INIT_RAM_13 = 256'h0E99AC528A300C032CC2588A0BAC200664422B0E0C2EBEA22EBA048891A4E384;
defparam prom_inst_2.INIT_RAM_14 = 256'h0C0370FFA2EBA66C0FF8B2AA2A9B23A912E321014581201C00402153ACA6372A;
defparam prom_inst_2.INIT_RAM_15 = 256'hB016D2F9690E4944081C16B090A6988088004A06F8CDB9BAE3B602622000C070;
defparam prom_inst_2.INIT_RAM_16 = 256'h2824A8E2EE38A28A2BA1CBB2ABE820688ACAD4E95460012845795AB8AAE9AE33;
defparam prom_inst_2.INIT_RAM_17 = 256'h3044AAAAAEBA418D052CCAB2AED658E3A0488862E1E3E2EEF0CE42AB332CB2CB;
defparam prom_inst_2.INIT_RAM_18 = 256'hA464ABB244A44AB90AEA0A85E17AAA00AE80A2AAABAEBA48E83C8DA22E929A02;
defparam prom_inst_2.INIT_RAM_19 = 256'hAD0A2AEC38EA223EB9F14F842ECEA123AECCEBBA223A44292E8BB3B39EAB1192;
defparam prom_inst_2.INIT_RAM_1A = 256'hAAD841692A4B91865AF07A20BBA0A01A8D0E804E18FBB4E86E1390A03B824408;
defparam prom_inst_2.INIT_RAM_1B = 256'h8528FAA38068806A8869101A26A492490A58962CC2AA288049882E88EE0A8840;
defparam prom_inst_2.INIT_RAM_1C = 256'h02996ACA9B1E5850B2FE1088EE492A91E0201A0680C0FA492A86184861B8DEAA;
defparam prom_inst_2.INIT_RAM_1D = 256'h723643EE20C99C1A287A54ECCBA4242A261622901A5896C2C8A69A499269B59A;
defparam prom_inst_2.INIT_RAM_1E = 256'hA1B2CCBC9A4A52BA7B1EC14CAE6A2E373882C1901198A28CC24B15A68292AEEB;
defparam prom_inst_2.INIT_RAM_1F = 256'hB88820861AEAAAABA0AE8AE81A62B22D1A21088AE2FEE8DA987B9B847B2E9808;
defparam prom_inst_2.INIT_RAM_20 = 256'h94949496208280C2492A86181C07082E9B41D1C92DE8924AAA861AEA112280B9;
defparam prom_inst_2.INIT_RAM_21 = 256'h08821A1A1A8187AB2EED91EC87B3984E350D0FCE88CC44AA223244AA72EAE8AA;
defparam prom_inst_2.INIT_RAM_22 = 256'h0A23F23C1ECCEE82FC8E330AA20B9080089682FBE8AA00001C1500C8BC228AA1;
defparam prom_inst_2.INIT_RAM_23 = 256'h9A8A44EE885A15872510F2F2FCDF3F2381AEE1CE23C5A2BC8AF0F2CCC0704AAA;
defparam prom_inst_2.INIT_RAM_24 = 256'h283AEBBB6E99BEDA061B7CB2CAA98A2BC52AA5A2A6882282A8A7882AF68BB873;
defparam prom_inst_2.INIT_RAM_25 = 256'hA4AD883A8A0A06062CC88409048416AF2F0F236CCAAAA21026D47C0ECCAF2F0F;
defparam prom_inst_2.INIT_RAM_26 = 256'h2AAC2492AA8A2AAEB633DC903AEAE380A3B0C77AE3678739ABA66D8067157AE2;
defparam prom_inst_2.INIT_RAM_27 = 256'h7EE2EFAA803BB4AF82D23CB210ECE43B308B81C80ADABAA3ACC2F23CA90BA832;
defparam prom_inst_2.INIT_RAM_28 = 256'hCE85BACEEE8EC072DEB8ACCCCECB8E2BD91C93E30893E948FA09CBE912ABA74A;
defparam prom_inst_2.INIT_RAM_29 = 256'hEA8EA8EACAB20A50B23A2A2B694BA3830E0C3830F2B3E3EA1EC87A3CC21A822C;
defparam prom_inst_2.INIT_RAM_2A = 256'h117E8AEC8784C4F0FA02A868687B33A32A32A32B33AEAAAFA182C3AF6AAB0B48;
defparam prom_inst_2.INIT_RAM_2B = 256'hB330BA3CBAB2BAEAEB9B2E6FBABAEA823AAC13F9F0033330B3B2500099233333;
defparam prom_inst_2.INIT_RAM_2C = 256'hB81825971A5FAACF303B333CCF33CB3251EEEECEECEECEE560341F36ADAB6ADB;
defparam prom_inst_2.INIT_RAM_2D = 256'hBEEC38A6F6188E18E18E2EFAEA2B2EAF2C3EC2EAD822BAFB0BC97B6D38A3CEB3;
defparam prom_inst_2.INIT_RAM_2E = 256'h8DA368B33A6632AAAC8F2033C8F23CB3308E8E8E81BCB00014BC72BB2BB2BA97;
defparam prom_inst_2.INIT_RAM_2F = 256'hA3CF38F2CCB30CC882B28A0A3E88FAE3AD372DCFAB34DB2EACD27CB3ACDA36B3;
defparam prom_inst_2.INIT_RAM_30 = 256'h48AA22304A86833B3A74AB328882EACE8728FB3A1E6CEB0C1EBAFCE063C580F5;
defparam prom_inst_2.INIT_RAM_31 = 256'hEEDA868E23ED8D8F6BA178AE86AB4AC8694EA13838383853B42E14E183C181D2;
defparam prom_inst_2.INIT_RAM_32 = 256'h8BC1AE330DA1EA2B3ADB68822DA88B7B707C8ECC9290D1EA842B8ACCECAD8D32;
defparam prom_inst_2.INIT_RAM_33 = 256'hA8CEA37688B0D38C34AE53220B2B8C0C9A2EB25AEA63613EBB95FAEE8EEB88CC;
defparam prom_inst_2.INIT_RAM_34 = 256'h34C120407BCAE80481AAB21BAA0E3F03FB522C1B0D2860DE8E4028B04B393A33;
defparam prom_inst_2.INIT_RAM_35 = 256'hC5E2C6CECB338E84B2E89BE1D991E89B61EE89B81EBFB8B603F81F62F0088812;
defparam prom_inst_2.INIT_RAM_36 = 256'hF6CCE0ABEEABACCBAB0BEEEEB2CAD366FC82FC96DB210AEA3E16EEBA801F1FC2;
defparam prom_inst_2.INIT_RAM_37 = 256'hEEEDBAEAE09B282CAC288AAEBBBAEAB3E267BE3ACDA70ABACC049EEEBB3853B3;
defparam prom_inst_2.INIT_RAM_38 = 256'h9350034040E0F09BAAC2F8ABA26FA0BAE3BBA1BAEEEA328FB213B2EECB0B6DBE;
defparam prom_inst_2.INIT_RAM_39 = 256'h2409BEEE0F2A212006BF337A7771B63CF2E06CBA842EBBBEE6102BA1390261E2;
defparam prom_inst_2.INIT_RAM_3A = 256'h8A6303802EBBAA2AA4A82800230D37B64E0200AE0800200AE00AE0000E243AEE;
defparam prom_inst_2.INIT_RAM_3B = 256'h9BBB87B52CC22424B3C8151A5AE78E00BAEEE00006680EB821B5515559858910;
defparam prom_inst_2.INIT_RAM_3C = 256'h106001104650002000698401920514004819081904200AEA802BAEE2DB8AECAA;
defparam prom_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFF0209044092FF901500EE46EE0146042FF8400049148;
defparam prom_inst_2.INIT_RAM_3E = 256'hFFFFE80FEF95AEEE91AA09B101FA6F6102DAD2D02D8B3050346DFB4E8F72D19E;
defparam prom_inst_2.INIT_RAM_3F = 256'hCCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hDF75D79F7DD75CCCFEEEECEDFFCEEEFE0FDFDDEDCCFDDCDDCDFECCEEEDFCFCDC;
defparam prom_inst_3.INIT_RAM_01 = 256'h565776575D57575755D5D7575757577575D55D57555DD7575D5D755D5D5D75E7;
defparam prom_inst_3.INIT_RAM_02 = 256'h555055555555552565565595D7595D7575D75D75D75D75D75D75D6ADD7AAD5D7;
defparam prom_inst_3.INIT_RAM_03 = 256'h8ACA9E8B2A728EEBA9AE8A6C1F848C3A30E82A08E8EC2FF85540050050554555;
defparam prom_inst_3.INIT_RAM_04 = 256'hD00EA5D0FAE3AB8F36F36F34524ACCAD9CE9EC33A624ACCAD2798847FBBAAFAA;
defparam prom_inst_3.INIT_RAM_05 = 256'h2A6A5A6AAAA32FDDFF661C947CA7A2B6D66652EA6A666A26C1B8D3DE0ABBC8EE;
defparam prom_inst_3.INIT_RAM_06 = 256'hC23227F7E7E3F33333E0B4F03F3999B166296FDB2D4D886666D32A0A666A6F2B;
defparam prom_inst_3.INIT_RAM_07 = 256'h8DCCC3082FA43BFECF32FFA62A23233A331473633262E56D64CD3FFFFFFF0D7F;
defparam prom_inst_3.INIT_RAM_08 = 256'hAAAE1859859B68BD3AAAA32B88E32B2F3AAA2667882C2BEB3ADFBF0BF7F26B71;
defparam prom_inst_3.INIT_RAM_09 = 256'h8CCCEBABD307A6222E3025BD08BB3330D3ECC9ED6ED616A2B8E4E59B0A66666A;
defparam prom_inst_3.INIT_RAM_0A = 256'hA691E7630C096863E386AFF23AF33ACFEA9CC4FFCD6EAABAA3ADB58CFC4A2D28;
defparam prom_inst_3.INIT_RAM_0B = 256'hFDF08F2EDABBAEDCE2C4CCF8AA8FBB069A6B4E3820ECCC3AB566EAA84AE38F29;
defparam prom_inst_3.INIT_RAM_0C = 256'hD52C8FFE1AAAAEEAD4E88F5D498BA96AAAAA8FB8C2D1AA898D825C9CA38F92B1;
defparam prom_inst_3.INIT_RAM_0D = 256'hE79A6971D4823BB8AEF78EB8E8B0662CBB488EB0D3DE0C69A69E7B02E74D4F5F;
defparam prom_inst_3.INIT_RAM_0E = 256'h98F88897CF42314EEECEDE3DE48CBC0EBCA3B338FF3FDFF99999898827CBB4B0;
defparam prom_inst_3.INIT_RAM_0F = 256'h4AAAAE28B1AA27A327A2BA8CAE8B53E0785BCAAAF3520C89480085885040B8D8;
defparam prom_inst_3.INIT_RAM_10 = 256'h992FFC2326F0BC22222FF38D08C4A2E34C4E1CDCDEDEDCCCE1AAEABAA2F2A8AB;
defparam prom_inst_3.INIT_RAM_11 = 256'hAA3673FF04F43322341082F74F3FC6BF2B8E3123FF23238ED73E131DE339D08C;
defparam prom_inst_3.INIT_RAM_12 = 256'h0423BB0F110CCEEAA22EEAAF2A9AAAB5F3CC432C08BCE3C2E0CD5EEAAE38B1AA;
defparam prom_inst_3.INIT_RAM_13 = 256'h4DAAB5FBC2EAFBAEDFB23BC35F0CCEE22AAEEF4CCCCD34E7CF38C87B98262336;
defparam prom_inst_3.INIT_RAM_14 = 256'h0A8230CBC2D34AAA0AC09BFFBFE723E2ABC32301551545500555455479E23A2C;
defparam prom_inst_3.INIT_RAM_15 = 256'h75356163AF48A6B910C8CAC328B8C0990BFCFB52E48100E3023CCCA1BDE0B82A;
defparam prom_inst_3.INIT_RAM_16 = 256'h965AE0DCDE15A69A6B8665D9B6AC7DAD1D9DB9B7FA2FF3E2577829C1E1B7651B;
defparam prom_inst_3.INIT_RAM_17 = 256'h24FC8820B8F312BC4EF9DAB6BC323BF78C87B8CFEDEFCDB4D488626AA69A69A6;
defparam prom_inst_3.INIT_RAM_18 = 256'hA545AF3865A65AF188EE48AFABE9F3569E19A6A78F38F0AC89314DAABCC54B52;
defparam prom_inst_3.INIT_RAM_19 = 256'h9F330BCF78D0B22EFBA2028FFEAEA223B2AAE2AAAAB8B62F6F0AAA128B8E5516;
defparam prom_inst_3.INIT_RAM_1A = 256'h5B1C9FFE1A27BE8EE8DCDEA89998B1334288A26E33ED3888B42218B12D0CA630;
defparam prom_inst_3.INIT_RAM_1B = 256'h8AE82B82029AACAA4466AB2A12ABAEBACAABAA266EABCAAC84AAA6AA6607A8CD;
defparam prom_inst_3.INIT_RAM_1C = 256'h520BA6BA4ACEE8EFA2373BAA66659F1BCCCC2A0A9090A9A69F1A698965B17F3B;
defparam prom_inst_3.INIT_RAM_1D = 256'hEEFEA3AB2A6C1F29AA69F76AAD2AEB16111422AFDAABAAA2A8B0F31FB26F3D8B;
defparam prom_inst_3.INIT_RAM_1E = 256'hA89AA6A66AA9AA6AE2388F7A96A9B4322BD752BB32BA6A7AA26ADDAAFAA2B62F;
defparam prom_inst_3.INIT_RAM_1F = 256'hB5C1E79A6BCAF38F1ABCF3CD4AFAF22F6AA98AEA7A30E0D9FBA96960A22A2888;
defparam prom_inst_3.INIT_RAM_20 = 256'h6B6B6B692E79C4CCA69E1A6BABEA79ED2B26AABAAE88A9A78F1A6BCE6AB068F2;
defparam prom_inst_3.INIT_RAM_21 = 256'hAAA22A2A2AD48DDB8AAE23AACAAA6A0CFDCDCEBEAAAA6626AAB0AAAA32E5D0B8;
defparam prom_inst_3.INIT_RAM_22 = 256'h8AABFC37376666A2FF0DD989AAA9A8AAAABD6AC21896AAAA2732B8AA4D556FD9;
defparam prom_inst_3.INIT_RAM_23 = 256'h4AAAAA66AA2B32B2B32B6E6CDB06FFCFB3B6726511BC2A5BA96C6266C4DCEEAA;
defparam prom_inst_3.INIT_RAM_24 = 256'h2F7CE2AB8E2AB4E3522928A9A78E1A6B1AEAEAAEBCAAAAA1AA9AA90AFA499C99;
defparam prom_inst_3.INIT_RAM_25 = 256'h689E09B8498D8DCDD666CAA44ECECC66E6D623C66AAE1B2A91FA9A4E666AEADA;
defparam prom_inst_3.INIT_RAM_26 = 256'h26CE2A6995A69F2AAAF6AC86F4E3C3332BB1DB34F789C994678AAE19AA2AF4F5;
defparam prom_inst_3.INIT_RAM_27 = 256'h8AE7CF387BAA989D0C62589B2E66539AABBBD3E0DAFAF38235E6623E198B8F78;
defparam prom_inst_3.INIT_RAM_28 = 256'hAAA23B3EAAAAE4F42D35AA9ADAD35EA7E248ABC330ABC48AF3D88BC48AAB0ABA;
defparam prom_inst_3.INIT_RAM_29 = 256'h9AA9AA9AA96A8BCC6AAAAAA8E88B02A30A8C2A30AA74A3BA48E06ACFA23AA21D;
defparam prom_inst_3.INIT_RAM_2A = 256'h202A8FF04A8888A89B526CECECEEB6AB6AB6AB6AB6999993B2A1DEB32222071A;
defparam prom_inst_3.INIT_RAM_2B = 256'h9998B47D3AB074EAD3AB4EAE3AB4EAAA5EB503E0482B0B098B1948024FD11113;
defparam prom_inst_3.INIT_RAM_2C = 256'hBD3A9000290E9AA6AA2AA69AA6A98999F695556966966960A8753C70AC2B0AC2;
defparam prom_inst_3.INIT_RAM_2D = 256'hE8882080DB20BA3BA3BA2EBBD2AC2E1F4F70A2EAE009FBD28B843B8D7D50DA6A;
defparam prom_inst_3.INIT_RAM_2E = 256'hA6A9A899B8AA32A29AA6AA29AA6A9899BDA6A6A6D4B128003DBDAAEAAEAAEACC;
defparam prom_inst_3.INIT_RAM_2F = 256'hBC96FB626667DAAAA236AA8AB848B8A3AC7F4E8FA6BFAA2E1AFEA8AA9A6A9A12;
defparam prom_inst_3.INIT_RAM_30 = 256'h889AAABD6AAA26AAB02BA6B8A898A9AD03EAC2BA08B1EBDD2A3B6B6CEDB3B863;
defparam prom_inst_3.INIT_RAM_31 = 256'h31E2C21F50AFBE0FEF803AB2B627DB08218893333B333B220DCCD88333A332CE;
defparam prom_inst_3.INIT_RAM_32 = 256'hCB53A2EA8E20822E74F0AAAAAD3A81B1B5B9A3348240D42188EB5AA9AF1E1E70;
defparam prom_inst_3.INIT_RAM_33 = 256'hAAE6AB92A8A8EC8E3B2A03AA8C2B48C04A2C34FBE3EF803F3880FCE2AEF3988E;
defparam prom_inst_3.INIT_RAM_34 = 256'h38C220A0878F0A09822AC203A2CCFCE3AACE8DAA8EC8ECE4BAAFC474AC0C2EB9;
defparam prom_inst_3.INIT_RAM_35 = 256'h4860694226B68E8970F0AB86E1A3F0AB40AD0ABD3A7C3AB803F40F0170248822;
defparam prom_inst_3.INIT_RAM_36 = 256'hB4AAF4AB4F2B4AA7468B4EEF34AACEAAA8933E46D382BAE2B825AF3B8084BD65;
defparam prom_inst_3.INIT_RAM_37 = 256'hAE6E34E6D4BBCAAAAA2AAAAD3ABCEAFB02E0B861527ECAB4AAC84AAF2AACEEAA;
defparam prom_inst_3.INIT_RAM_38 = 256'h2BC801C6C6C5E4AB46A2C0ABC2AF18B4D79BC074E6F1B582B406B4E6D28B4E38;
defparam prom_inst_3.INIT_RAM_39 = 256'h6767C33CC8F6F3F0269651935297169311F41D398ADD3AB8EA2B6BC06B1B6909;
defparam prom_inst_3.INIT_RAM_3A = 256'h88EB723BB0E3999B422A26489AAFEBE2222622E62A22622EA22EE2222E2ABB8E;
defparam prom_inst_3.INIT_RAM_3B = 256'hC199CDDA26622210F78CB8CBCB4388EEC38E6AAAA22C4ED0C3F320CCA8CCC888;
defparam prom_inst_3.INIT_RAM_3C = 256'h554555515455500555411555145554015151515154122E6D08BAB8EAD1EA72B4;
defparam prom_inst_3.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFF0051555514001555500054005554554001500551550;
defparam prom_inst_3.INIT_RAM_3E = 256'hFFFFD401551515451515444332C113E330F9F9F30F9D71F737CEC3FC0F62FAAE;
defparam prom_inst_3.INIT_RAM_3F = 256'hCCCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

endmodule //basicRom
